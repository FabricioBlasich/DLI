library ieee;
use ieee.std_logic_1164.all;


entity Ejercicio_Lab2 is

	generic
	(
		DATA_WIDTH : natural := 8
	);

	port 
	(

	);

end entity;

architecture a_Ejercicio_Lab2 of Ejercicio_Lab2 is

component deco
	A, B, C, D	   : in std_logic;
	

end component;
begin
end Ejercicio_Lab2;
